--==============================================================================
--== Logisim-evolution goes FPGA automatic generated VHDL code                ==
--== https://github.com/logisim-evolution/                                    ==
--==                                                                          ==
--==                                                                          ==
--== Project   : print_ADXL345_values                                         ==
--== Component : random_tb                                                    ==
--==                                                                          ==
--==============================================================================


LIBRARY ieee;
USE ieee.std_logic_1164.all;
USE ieee.numeric_std.all;


ENTITY random_tb IS
   PORT ( Input_1      : IN  std_logic;
          Output_bus_1 : OUT std_logic_vector( 7 DOWNTO 0 ) );
END ENTITY random_tb;
