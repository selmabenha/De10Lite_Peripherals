--==============================================================================
--== Logisim-evolution goes FPGA automatic generated VHDL code                ==
--== https://github.com/logisim-evolution/                                    ==
--==                                                                          ==
--==                                                                          ==
--== Project   : get_to_zero                                                  ==
--== Component : logisimTopLevelShell                                         ==
--==                                                                          ==
--==============================================================================


LIBRARY ieee;
USE ieee.std_logic_1164.all;
USE ieee.numeric_std.all;


ENTITY logisimTopLevelShell IS
   PORT ( enable_0                                  : IN  std_logic;
          fpgaGlobalClock                           : IN  std_logic;
          reset_0                                   : IN  std_logic;
          stop_0                                    : IN  std_logic;
          n_hex0_L_7_Segment_Display_1_DecimalPoint : OUT std_logic;
          n_hex0_L_7_Segment_Display_1_Segment_A    : OUT std_logic;
          n_hex0_L_7_Segment_Display_1_Segment_B    : OUT std_logic;
          n_hex0_L_7_Segment_Display_1_Segment_C    : OUT std_logic;
          n_hex0_L_7_Segment_Display_1_Segment_D    : OUT std_logic;
          n_hex0_L_7_Segment_Display_1_Segment_E    : OUT std_logic;
          n_hex0_L_7_Segment_Display_1_Segment_F    : OUT std_logic;
          n_hex0_L_7_Segment_Display_1_Segment_G    : OUT std_logic;
          n_hex1_L_7_Segment_Display_1_DecimalPoint : OUT std_logic;
          n_hex1_L_7_Segment_Display_1_Segment_A    : OUT std_logic;
          n_hex1_L_7_Segment_Display_1_Segment_B    : OUT std_logic;
          n_hex1_L_7_Segment_Display_1_Segment_C    : OUT std_logic;
          n_hex1_L_7_Segment_Display_1_Segment_D    : OUT std_logic;
          n_hex1_L_7_Segment_Display_1_Segment_E    : OUT std_logic;
          n_hex1_L_7_Segment_Display_1_Segment_F    : OUT std_logic;
          n_hex1_L_7_Segment_Display_1_Segment_G    : OUT std_logic;
          n_hex2_L_7_Segment_Display_1_DecimalPoint : OUT std_logic;
          n_hex2_L_7_Segment_Display_1_Segment_A    : OUT std_logic;
          n_hex2_L_7_Segment_Display_1_Segment_B    : OUT std_logic;
          n_hex2_L_7_Segment_Display_1_Segment_C    : OUT std_logic;
          n_hex2_L_7_Segment_Display_1_Segment_D    : OUT std_logic;
          n_hex2_L_7_Segment_Display_1_Segment_E    : OUT std_logic;
          n_hex2_L_7_Segment_Display_1_Segment_F    : OUT std_logic;
          n_hex2_L_7_Segment_Display_1_Segment_G    : OUT std_logic );
END ENTITY logisimTopLevelShell;
