--==============================================================================
--== Logisim-evolution goes FPGA automatic generated VHDL code                ==
--== https://github.com/logisim-evolution/                                    ==
--==                                                                          ==
--==                                                                          ==
--== Project   : get_to_zero                                                  ==
--== Component : counter_fsm                                                  ==
--==                                                                          ==
--==============================================================================


LIBRARY ieee;
USE ieee.std_logic_1164.all;
USE ieee.numeric_std.all;


ENTITY counter_fsm IS
   PORT ( logisimClockTree0 : IN  std_logic_vector( 4 DOWNTO 0 );
          reset             : IN  std_logic;
          state_1           : IN  std_logic;
          state_2           : IN  std_logic;
          state_3           : IN  std_logic;
          state_output      : OUT std_logic_vector( 1 DOWNTO 0 ) );
END ENTITY counter_fsm;
