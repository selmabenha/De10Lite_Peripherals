--==============================================================================
--== Logisim-evolution goes FPGA automatic generated VHDL code                ==
--== https://github.com/logisim-evolution/                                    ==
--==                                                                          ==
--==                                                                          ==
--== Project   : accelerometer_v2                                             ==
--== Component : sevenseg_numbers_logic                                       ==
--==                                                                          ==
--==============================================================================


LIBRARY ieee;
USE ieee.std_logic_1164.all;
USE ieee.numeric_std.all;


ENTITY sevenseg_numbers_logic IS
   PORT ( accel        : IN  std_logic_vector( 3 DOWNTO 0 );
          sevensegment : OUT std_logic_vector( 7 DOWNTO 0 ) );
END ENTITY sevenseg_numbers_logic;
