--==============================================================================
--== Logisim-evolution goes FPGA automatic generated VHDL code                ==
--== https://github.com/logisim-evolution/                                    ==
--==                                                                          ==
--==                                                                          ==
--== Project   : Inshallah                                                    ==
--== Component : logisimTopLevelShell                                         ==
--==                                                                          ==
--==============================================================================


LIBRARY ieee;
USE ieee.std_logic_1164.all;
USE ieee.numeric_std.all;


ENTITY logisimTopLevelShell IS
   PORT ( fpgaGlobalClock  : IN  std_logic;
          n_Input_bus_1_0  : IN  std_logic;
          n_Input_bus_1_1  : IN  std_logic;
          n_Output_bus_1_0 : OUT std_logic;
          n_Output_bus_1_1 : OUT std_logic;
          n_Output_bus_1_2 : OUT std_logic;
          n_Output_bus_1_3 : OUT std_logic;
          n_Output_bus_1_4 : OUT std_logic;
          n_Output_bus_1_5 : OUT std_logic;
          n_Output_bus_1_6 : OUT std_logic;
          n_Output_bus_1_7 : OUT std_logic );
END ENTITY logisimTopLevelShell;
