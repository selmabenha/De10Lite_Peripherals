--==============================================================================
--== Logisim-evolution goes FPGA automatic generated VHDL code                ==
--== https://github.com/logisim-evolution/                                    ==
--==                                                                          ==
--==                                                                          ==
--== Project   : division                                                     ==
--== Component : memory_test                                                  ==
--==                                                                          ==
--==============================================================================


LIBRARY ieee;
USE ieee.std_logic_1164.all;
USE ieee.numeric_std.all;


ENTITY memory_test IS
   PORT ( Input_1  : IN  std_logic;
          Input_2  : IN  std_logic;
          Output_1 : OUT std_logic );
END ENTITY memory_test;
